module CMOSCamera( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  output       io_lcdSpi_serialClock, // @[:@6.4]
  output       io_lcdSpi_dataCommand, // @[:@6.4]
  output       io_lcdSpi_chipSelectN, // @[:@6.4]
  output       io_lcdSpi_masterOutSlaveIn, // @[:@6.4]
  input        io_lcdSpi_masterInSlaveOut, // @[:@6.4]
  output       io_lcdSpi_resetN, // @[:@6.4]
  output       io_lcdSpi_backLight, // @[:@6.4]
  output       io_cmosCam_systemClock, // @[:@6.4]
  input        io_cmosCam_verticalSync, // @[:@6.4]
  input        io_cmosCam_horizontalRef, // @[:@6.4]
  input        io_cmosCam_pixelclock, // @[:@6.4]
  input  [7:0] io_cmosCam_pixcelData, // @[:@6.4]
  output       io_cmosCam_sccbClock, // @[:@6.4]
  output       io_cmosCam_sccbData, // @[:@6.4]
  output       io_cmosCam_resetN, // @[:@6.4]
  output       io_cmosCam_powerDown // @[:@6.4]
);
  assign io_lcdSpi_serialClock = 1'h1; // @[CMOSCamera.scala 36:25:@8.4]
  assign io_lcdSpi_dataCommand = 1'h1; // @[CMOSCamera.scala 37:25:@9.4]
  assign io_lcdSpi_chipSelectN = 1'h1; // @[CMOSCamera.scala 38:25:@10.4]
  assign io_lcdSpi_masterOutSlaveIn = 1'h1; // @[CMOSCamera.scala 39:30:@11.4]
  assign io_lcdSpi_resetN = 1'h1; // @[CMOSCamera.scala 40:20:@12.4]
  assign io_lcdSpi_backLight = 1'h1; // @[CMOSCamera.scala 41:23:@13.4]
  assign io_cmosCam_systemClock = 1'h1; // @[CMOSCamera.scala 43:26:@14.4]
  assign io_cmosCam_sccbClock = 1'h1; // @[CMOSCamera.scala 44:24:@15.4]
  assign io_cmosCam_sccbData = 1'h1; // @[CMOSCamera.scala 45:23:@16.4]
  assign io_cmosCam_resetN = 1'h1; // @[CMOSCamera.scala 46:21:@17.4]
  assign io_cmosCam_powerDown = 1'h0; // @[CMOSCamera.scala 47:24:@18.4]
endmodule
